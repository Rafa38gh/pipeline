-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.


-- Generated by Quartus Prime Version 20.1 (Build Build 720 11/11/2020)
-- Created on Fri Nov 21 10:37:39 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE full_adder_package IS
	COMPONENT full_adder
		PORT
		(
			CIN		:	 IN STD_LOGIC;
			X		:	 IN STD_LOGIC;
			Y		:	 IN STD_LOGIC;
			COUT		:	 OUT STD_LOGIC;
			S		:	 OUT STD_LOGIC
		);
	END COMPONENT;
END PACKAGE;