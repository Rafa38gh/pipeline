-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.


-- Generated by Quartus Prime Version 20.1 (Build Build 720 11/11/2020)
-- Created on Fri Nov 21 15:10:19 2025
LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE UC_package IS
	COMPONENT UC
		PORT
		(
			OPCODE		:	 IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			REGDST		:	 OUT STD_LOGIC;
			REGWRITE		:	 OUT STD_LOGIC;
			MEMREAD		:	 OUT STD_LOGIC;
			MEMWRITE		:	 OUT STD_LOGIC;
			MEMTOREG		:	 OUT STD_LOGIC;
			BRANCH		:	 OUT STD_LOGIC;
			JUMP		:	 OUT STD_LOGIC;
			ALUSRC		:	 OUT STD_LOGIC;
			ALUOP			:	 OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
		);
	END COMPONENT;
END PACKAGE;