-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.


-- Generated by Quartus Prime Version 20.1 (Build Build 720 11/11/2020)
-- Created on Mon Dec 01 12:23:31 2025
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;
USE work.pc_package.all;
USE work.mem_inst_package.all;
USE work.ULA_sim_package.all;
USE work.pipe_reg_package.all;
USE work.reg_file_package.all;
USE work.UC_package.all;
USE work.mux2_1_package.all;
USE work.ULA16_package.all;
USE work.data_mem_package.all;

PACKAGE pipeline_package IS
	COMPONENT pipeline
		PORT
		(
			CLK		:	 IN STD_LOGIC;
			RESET		:	 IN STD_LOGIC;
			ENABLE		:	 IN STD_LOGIC;
			RS		:	 OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
			RT		:	 OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
		);
	END COMPONENT;
END PACKAGE;